/** @module : phi
 *  @author : Secure Trusted and Assured Microelectronics (STAM) Center

 *  Copyright (c) 2023 PQC.Secure (STAM/SCAI/ASU)
 *  Permission is hereby granted, free of charge, to any person obtaining a copy
 *  of this software and associated documentation files (the "Software"), to deal
 *  in the Software without restriction, including without limitation the rights
 *  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 *  copies of the Software, and to permit persons to whom the Software is
 *  furnished to do so, subject to the following conditions:
 *  The above copyright notice and this permission notice shall be included in
 *  all copies or substantial portions of the Software.
 z
 *  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 *  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 *  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 *  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 *  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 *  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 *  THE SOFTWARE.
 *
 *
 */

/*********************************************************************************
*                                         phi                                    *
*********************************************************************************/



// for 2*N = 16, p = 17
if (N == 8)
begin
    // phi = 3 for 2*N = 16, p = 17
    phi[0] <= 1; phi[1] <= 3; phi[2] <= 9; phi[3] <= 10; phi[4] <= 13; phi[5] <= 5; phi[6] <= 15; phi[7] <= 11;
    // phi[16] == 1
    
    
    // iphi = 6 for 2*N = 16, p = 17
    iphi[0] <= 1; iphi[1] <= 6; iphi[2] <= 2; iphi[3] <= 12; iphi[4] <= 4; iphi[5] <= 7; iphi[6] <= 8; iphi[7] <= 14;
    // iphi[16] == 1
end


// for 2*N = 32, p = 97
else if (N == 16)
begin
    // phi = 28 for 2*N = 32, p = 97
    phi[0] <= 1; phi[1] <= 28; phi[2] <= 8; phi[3] <= 30; phi[4] <= 64; phi[5] <= 46; phi[6] <= 27; phi[7] <= 77; 
    phi[8] <= 22; phi[9] <= 34; phi[10] <= 79; phi[11] <= 78; phi[12] <= 50; phi[13] <= 42; phi[14] <= 12; phi[15] <= 45;
    // phi[32] == 1
    
    // phi = 52 for 2*N = 32, p = 97
    iphi[0] <= 1; iphi[1] <= 52; iphi[2] <= 85; iphi[3] <= 55; iphi[4] <= 47; iphi[5] <= 19; iphi[6] <= 18; iphi[7] <= 63; 
    iphi[8] <= 75; iphi[9] <= 20; iphi[10] <= 70; iphi[11] <= 51; iphi[12] <= 33; iphi[13] <= 67; iphi[14] <= 89; iphi[15] <= 69;
    // iphi[32] == 1
end


// for 2*N = 64, p = 193
else if (N == 32)
begin
    phi[0] <= 1; phi[1] <= 125; phi[2] <= 185; phi[3] <= 158; phi[4] <= 64; phi[5] <= 87; phi[6] <= 67; phi[7] <= 76; 
    phi[8] <= 43; phi[9] <= 164; phi[10] <= 42; phi[11] <= 39; phi[12] <= 50; phi[13] <= 74; phi[14] <= 179; phi[15] <= 180; 
    phi[16] <= 112; phi[17] <= 104; phi[18] <= 69; phi[19] <= 133; phi[20] <= 27; phi[21] <= 94; phi[22] <= 170; phi[23] <= 20; 
    phi[24] <= 184; phi[25] <= 33; phi[26] <= 72; phi[27] <= 122; phi[28] <= 3; phi[29] <= 182; phi[30] <= 169; phi[31] <= 88;
    
    iphi[0] <= 1; iphi[1] <= 105; iphi[2] <= 24; iphi[3] <= 11; iphi[4] <= 190; iphi[5] <= 71; iphi[6] <= 121; iphi[7] <= 160; 
    iphi[8] <= 9; iphi[9] <= 173; iphi[10] <= 23; iphi[11] <= 99; iphi[12] <= 166; iphi[13] <= 60; iphi[14] <= 124; iphi[15] <= 89; 
    iphi[16] <= 81; iphi[17] <= 13; iphi[18] <= 14; iphi[19] <= 119; iphi[20] <= 143; iphi[21] <= 154; iphi[22] <= 151; iphi[23] <= 29; 
    iphi[24] <= 150; iphi[25] <= 117; iphi[26] <= 126; iphi[27] <= 106; iphi[28] <= 129; iphi[29] <= 35; iphi[30] <= 8; iphi[31] <= 68;
end


// for 2*N = 128, 
else if (N == 64)
begin
    // p = 257
    /*
    phi[0] <= 1; phi[1] <= 9; phi[2] <= 81; phi[3] <= 215; phi[4] <= 136; phi[5] <= 196; phi[6] <= 222; phi[7] <= 199; 
    phi[8] <= 249; phi[9] <= 185; phi[10] <= 123; phi[11] <= 79; phi[12] <= 197; phi[13] <= 231; phi[14] <= 23; phi[15] <= 207; 
    phi[16] <= 64; phi[17] <= 62; phi[18] <= 44; phi[19] <= 139; phi[20] <= 223; phi[21] <= 208; phi[22] <= 73; phi[23] <= 143; 
    phi[24] <= 2; phi[25] <= 18; phi[26] <= 162; phi[27] <= 173; phi[28] <= 15; phi[29] <= 135; phi[30] <= 187; phi[31] <= 141; 
    phi[32] <= 241; phi[33] <= 113; phi[34] <= 246; phi[35] <= 158; phi[36] <= 137; phi[37] <= 205; phi[38] <= 46; phi[39] <= 157; 
    phi[40] <= 128; phi[41] <= 124; phi[42] <= 88; phi[43] <= 21; phi[44] <= 189; phi[45] <= 159; phi[46] <= 146; phi[47] <= 29; 
    phi[48] <= 4; phi[49] <= 36; phi[50] <= 67; phi[51] <= 89; phi[52] <= 30; phi[53] <= 13; phi[54] <= 117; phi[55] <= 25; 
    phi[56] <= 225; phi[57] <= 226; phi[58] <= 235; phi[59] <= 59; phi[60] <= 17; phi[61] <= 153; phi[62] <= 92; phi[63] <= 57;
    
    iphi[0] <= 1; iphi[1] <= 200; iphi[2] <= 165; iphi[3] <= 104; iphi[4] <= 240; iphi[5] <= 198; iphi[6] <= 22; iphi[7] <= 31; 
    iphi[8] <= 32; iphi[9] <= 232; iphi[10] <= 140; iphi[11] <= 244; iphi[12] <= 227; iphi[13] <= 168; iphi[14] <= 190; iphi[15] <= 221; 
    iphi[16] <= 253; iphi[17] <= 228; iphi[18] <= 111; iphi[19] <= 98; iphi[20] <= 68; iphi[21] <= 236; iphi[22] <= 169; iphi[23] <= 133; 
    iphi[24] <= 129; iphi[25] <= 100; iphi[26] <= 211; iphi[27] <= 52; iphi[28] <= 120; iphi[29] <= 99; iphi[30] <= 11; iphi[31] <= 144; 
    iphi[32] <= 16; iphi[33] <= 116; iphi[34] <= 70; iphi[35] <= 122; iphi[36] <= 242; iphi[37] <= 84; iphi[38] <= 95; iphi[39] <= 239; 
    iphi[40] <= 255; iphi[41] <= 114; iphi[42] <= 184; iphi[43] <= 49; iphi[44] <= 34; iphi[45] <= 118; iphi[46] <= 213; iphi[47] <= 195; 
    iphi[48] <= 193; iphi[49] <= 50; iphi[50] <= 234; iphi[51] <= 26; iphi[52] <= 60; iphi[53] <= 178; iphi[54] <= 134; iphi[55] <= 72; 
    iphi[56] <= 8; iphi[57] <= 58; iphi[58] <= 35; iphi[59] <= 61; iphi[60] <= 121; iphi[61] <= 42; iphi[62] <= 176; iphi[63] <= 248;
    */
    
    // p == 1153
    phi[0] <= 1; phi[1] <= 1096; phi[2] <= 943; phi[3] <= 440; phi[4] <= 286; phi[5] <= 993; phi[6] <= 1049; phi[7] <= 163; 
    phi[8] <= 1086; phi[9] <= 360; phi[10] <= 234; phi[11] <= 498; phi[12] <= 439; phi[13] <= 343; phi[14] <= 50; phi[15] <= 609; 
    phi[16] <= 1030; phi[17] <= 93; phi[18] <= 464; phi[19] <= 71; phi[20] <= 565; phi[21] <= 79; phi[22] <= 109; phi[23] <= 705; 
    phi[24] <= 170; phi[25] <= 687; phi[26] <= 43; phi[27] <= 1008; phi[28] <= 194; phi[29] <= 472; phi[30] <= 768; phi[31] <= 38; 
    phi[32] <= 140; phi[33] <= 91; phi[34] <= 578; phi[35] <= 491; phi[36] <= 838; phi[37] <= 660; phi[38] <= 429; phi[39] <= 913;
    phi[40] <= 997; phi[41] <= 821; phi[42] <= 476; phi[43] <= 540; phi[44] <= 351; phi[45] <= 747; phi[46] <= 82; phi[47] <= 1091; 
    phi[48] <= 75; phi[49] <= 337; phi[50] <= 392; phi[51] <= 716; phi[52] <= 696; phi[53] <= 683; phi[54] <= 271; phi[55] <= 695; 
    phi[56] <= 740; phi[57] <= 481; phi[58] <= 255; phi[59] <= 454; phi[60] <= 641; phi[61] <= 359; phi[62] <= 291; phi[63] <= 708;
     
    iphi[0] <= 1; iphi[1] <= 445; iphi[2] <= 862; iphi[3] <= 794; iphi[4] <= 512; iphi[5] <= 699; iphi[6] <= 898; iphi[7] <= 672; 
    iphi[8] <= 413; iphi[9] <= 458; iphi[10] <= 882; iphi[11] <= 470; iphi[12] <= 457; iphi[13] <= 437; iphi[14] <= 761; iphi[15] <= 816; 
    iphi[16] <= 1078; iphi[17] <= 62; iphi[18] <= 1071; iphi[19] <= 406; iphi[20] <= 802; iphi[21] <= 613; iphi[22] <= 677; iphi[23] <= 332; 
    iphi[24] <= 156; iphi[25] <= 240; iphi[26] <= 724; iphi[27] <= 493; iphi[28] <= 315; iphi[29] <= 662; iphi[30] <= 575; iphi[31] <= 1062; 
    iphi[32] <= 1013; iphi[33] <= 1115; iphi[34] <= 385; iphi[35] <= 681; iphi[36] <= 959; iphi[37] <= 145; iphi[38] <= 1110; iphi[39] <= 466; 
    iphi[40] <= 983; iphi[41] <= 448; iphi[42] <= 1044; iphi[43] <= 1074; iphi[44] <= 588; iphi[45] <= 1082; iphi[46] <= 689; iphi[47] <= 1060; 
    iphi[48] <= 123; iphi[49] <= 544; iphi[50] <= 1103; iphi[51] <= 810; iphi[52] <= 714; iphi[53] <= 655; iphi[54] <= 919; iphi[55] <= 793; 
    iphi[56] <= 67; iphi[57] <= 990; iphi[58] <= 104; iphi[59] <= 160; iphi[60] <= 867; iphi[61] <= 713; iphi[62] <= 210; iphi[63] <= 57;
end



// for 2*N = 256, p = 769
else if (N == 128)
begin
    if (p == 769)
    begin
        phi[0] <= 1; phi[1] <= 343; phi[2] <= 761; phi[3] <= 332; phi[4] <= 64; phi[5] <= 420; phi[6] <= 257; phi[7] <= 485; 
        phi[8] <= 251; phi[9] <= 734; phi[10] <= 299; phi[11] <= 280; phi[12] <= 684; phi[13] <= 67; phi[14] <= 680; phi[15] <= 233; 
        phi[16] <= 712; phi[17] <= 443; phi[18] <= 456; phi[19] <= 301; phi[20] <= 197; phi[21] <= 668; phi[22] <= 731; phi[23] <= 39; 
        phi[24] <= 304; phi[25] <= 457; phi[26] <= 644; phi[27] <= 189; phi[28] <= 231; phi[29] <= 26; phi[30] <= 459; phi[31] <= 561; 
        phi[32] <= 173; phi[33] <= 126; phi[34] <= 154; phi[35] <= 530; phi[36] <= 306; phi[37] <= 374; phi[38] <= 628; phi[39] <= 84; 
        phi[40] <= 359; phi[41] <= 97; phi[42] <= 204; phi[43] <= 762; phi[44] <= 675; phi[45] <= 56; phi[46] <= 752; phi[47] <= 321; 
        phi[48] <= 136; phi[49] <= 508; phi[50] <= 450; phi[51] <= 550; phi[52] <= 245; phi[53] <= 214; phi[54] <= 347; phi[55] <= 595; 
        phi[56] <= 300; phi[57] <= 623; phi[58] <= 676; phi[59] <= 399; phi[60] <= 744; phi[61] <= 653; phi[62] <= 200; phi[63] <= 159; 
        phi[64] <= 707; phi[65] <= 266; phi[66] <= 496; phi[67] <= 179; phi[68] <= 646; phi[69] <= 106; phi[70] <= 215; phi[71] <= 690; 
        phi[72] <= 587; phi[73] <= 632; phi[74] <= 687; phi[75] <= 327; phi[76] <= 656; phi[77] <= 460; phi[78] <= 135; phi[79] <= 165; 
        phi[80] <= 458; phi[81] <= 218; phi[82] <= 181; phi[83] <= 563; phi[84] <= 90; phi[85] <= 110; phi[86] <= 49; phi[87] <= 658; 
        phi[88] <= 377; phi[89] <= 119; phi[90] <= 60; phi[91] <= 586; phi[92] <= 289; phi[93] <= 695; phi[94] <= 764; phi[95] <= 592; 
        phi[96] <= 40; phi[97] <= 647; phi[98] <= 449; phi[99] <= 207; phi[100] <= 253; phi[101] <= 651; phi[102] <= 283; phi[103] <= 175; 
        phi[104] <= 43; phi[105] <= 138; phi[106] <= 425; phi[107] <= 434; phi[108] <= 445; phi[109] <= 373; phi[110] <= 285; phi[111] <= 92; 
        phi[112] <= 27; phi[113] <= 33; phi[114] <= 553; phi[115] <= 505; phi[116] <= 190; phi[117] <= 574; phi[118] <= 18; phi[119] <= 22; 
        phi[120] <= 625; phi[121] <= 593; phi[122] <= 383; phi[123] <= 639; phi[124] <= 12; phi[125] <= 271; phi[126] <= 673; phi[127] <= 139;
        
        iphi[0] <= 1; iphi[1] <= 630; iphi[2] <= 96; iphi[3] <= 498; iphi[4] <= 757; iphi[5] <= 130; iphi[6] <= 386; iphi[7] <= 176; 
        iphi[8] <= 144; iphi[9] <= 747; iphi[10] <= 751; iphi[11] <= 195; iphi[12] <= 579; iphi[13] <= 264; iphi[14] <= 216; iphi[15] <= 736; 
        iphi[16] <= 742; iphi[17] <= 677; iphi[18] <= 484; iphi[19] <= 396; iphi[20] <= 324; iphi[21] <= 335; iphi[22] <= 344; iphi[23] <= 631; 
        iphi[24] <= 726; iphi[25] <= 594; iphi[26] <= 486; iphi[27] <= 118; iphi[28] <= 516; iphi[29] <= 562; iphi[30] <= 320; iphi[31] <= 122; 
        iphi[32] <= 729; iphi[33] <= 177; iphi[34] <= 5; iphi[35] <= 74; iphi[36] <= 480; iphi[37] <= 183; iphi[38] <= 709; iphi[39] <= 650; 
        iphi[40] <= 392; iphi[41] <= 111; iphi[42] <= 720; iphi[43] <= 659; iphi[44] <= 679; iphi[45] <= 206; iphi[46] <= 588; iphi[47] <= 551; 
        iphi[48] <= 311; iphi[49] <= 604; iphi[50] <= 634; iphi[51] <= 309; iphi[52] <= 113; iphi[53] <= 442; iphi[54] <= 82; iphi[55] <= 137; 
        iphi[56] <= 182; iphi[57] <= 79; iphi[58] <= 554; iphi[59] <= 663; iphi[60] <= 123; iphi[61] <= 590; iphi[62] <= 273; iphi[63] <= 503; 
        iphi[64] <= 62; iphi[65] <= 610; iphi[66] <= 569; iphi[67] <= 116; iphi[68] <= 25; iphi[69] <= 370; iphi[70] <= 93; iphi[71] <= 146; 
        iphi[72] <= 469; iphi[73] <= 174; iphi[74] <= 422; iphi[75] <= 555; iphi[76] <= 524; iphi[77] <= 219; iphi[78] <= 319; iphi[79] <= 261; 
        iphi[80] <= 633; iphi[81] <= 448; iphi[82] <= 17; iphi[83] <= 713; iphi[84] <= 94; iphi[85] <= 7; iphi[86] <= 565; iphi[87] <= 672; 
        iphi[88] <= 410; iphi[89] <= 685; iphi[90] <= 141; iphi[91] <= 395; iphi[92] <= 463; iphi[93] <= 239; iphi[94] <= 615; iphi[95] <= 643; 
        iphi[96] <= 596; iphi[97] <= 208; iphi[98] <= 310; iphi[99] <= 743; iphi[100] <= 538; iphi[101] <= 580; iphi[102] <= 125; iphi[103] <= 312; 
        iphi[104] <= 465; iphi[105] <= 730; iphi[106] <= 38; iphi[107] <= 101; iphi[108] <= 572; iphi[109] <= 468; iphi[110] <= 313; iphi[111] <= 326; 
        iphi[112] <= 57; iphi[113] <= 536; iphi[114] <= 89; iphi[115] <= 702; iphi[116] <= 85; iphi[117] <= 489; iphi[118] <= 470; iphi[119] <= 35; 
        iphi[120] <= 518; iphi[121] <= 284; iphi[122] <= 512; iphi[123] <= 349; iphi[124] <= 705; iphi[125] <= 437; iphi[126] <= 8; iphi[127] <= 426;
    end
    
    else if (p == 3329)
    begin
        phi[0] <= 1; phi[1] <= 3061; phi[2] <= 1915; phi[3] <= 2775; phi[4] <= 1996; phi[5] <= 1041; phi[6] <= 648; phi[7] <= 2773; 
        phi[8] <= 2532; phi[9] <= 540; phi[10] <= 1756; phi[11] <= 2110; phi[12] <= 450; phi[13] <= 2573; phi[14] <= 2868; phi[15] <= 375; 
        phi[16] <= 2699; phi[17] <= 2390; phi[18] <= 1977; phi[19] <= 2804; phi[20] <= 882; phi[21] <= 3312; phi[22] <= 1227; phi[23] <= 735; 
        phi[24] <= 2760; phi[25] <= 2687; phi[26] <= 2277; phi[27] <= 2300; phi[28] <= 2794; phi[29] <= 233; phi[30] <= 807; phi[31] <= 109; 
        phi[32] <= 749; phi[33] <= 2337; phi[34] <= 2865; phi[35] <= 1179; phi[36] <= 283; phi[37] <= 723; phi[38] <= 2647; phi[39] <= 3010; 
        phi[40] <= 2267; phi[41] <= 1651; phi[42] <= 289; phi[43] <= 2444; phi[44] <= 821; phi[45] <= 3015; phi[46] <= 927; phi[47] <= 1239; 
        phi[48] <= 848; phi[49] <= 2437; phi[50] <= 2697; phi[51] <= 2926; phi[52] <= 1476; phi[53] <= 583; phi[54] <= 219; phi[55] <= 1230; 
        phi[56] <= 3260; phi[57] <= 1847; phi[58] <= 1025; phi[59] <= 1607; phi[60] <= 2094; phi[61] <= 1409; phi[62] <= 1894; phi[63] <= 1745; 
        phi[64] <= 1729; phi[65] <= 2688; phi[66] <= 2009; phi[67] <= 886; phi[68] <= 2240; phi[69] <= 2229; phi[70] <= 1848; phi[71] <= 757; 
        phi[72] <= 193; phi[73] <= 1540; phi[74] <= 76; phi[75] <= 2935; phi[76] <= 2393; phi[77] <= 1173; phi[78] <= 1891; phi[79] <= 2549; 
        phi[80] <= 2642; phi[81] <= 1021; phi[82] <= 2679; phi[83] <= 1092; phi[84] <= 296; phi[85] <= 568; phi[86] <= 910; phi[87] <= 2466; 
        phi[88] <= 1583; phi[89] <= 1868; phi[90] <= 2055; phi[91] <= 1874; phi[92] <= 447; phi[93] <= 48; phi[94] <= 452; phi[95] <= 2037; 
        phi[96] <= 40; phi[97] <= 2596; phi[98] <= 33; phi[99] <= 1143; phi[100] <= 3273; phi[101] <= 1692; phi[102] <= 2617; phi[103] <= 1063; 
        phi[104] <= 1410; phi[105] <= 1626; phi[106] <= 331; phi[107] <= 1175; phi[108] <= 1355; phi[109] <= 3050; phi[110] <= 1534; phi[111] <= 1684; 
        phi[112] <= 1432; phi[113] <= 2388; phi[114] <= 2513; phi[115] <= 2303; phi[116] <= 1990; phi[117] <= 2649; phi[118] <= 2474; phi[119] <= 2768; 
        phi[120] <= 543; phi[121] <= 952; phi[122] <= 1197; phi[123] <= 2117; phi[124] <= 1903; phi[125] <= 2662; phi[126] <= 2319; phi[127] <= 1031;
        
        iphi[0] <= 1; iphi[1] <= 2298; iphi[2] <= 1010; iphi[3] <= 667; iphi[4] <= 1426; iphi[5] <= 1212; iphi[6] <= 2132; iphi[7] <= 2377; 
        iphi[8] <= 2786; iphi[9] <= 561; iphi[10] <= 855; iphi[11] <= 680; iphi[12] <= 1339; iphi[13] <= 1026; iphi[14] <= 816; iphi[15] <= 941; 
        iphi[16] <= 1897; iphi[17] <= 1645; iphi[18] <= 1795; iphi[19] <= 279; iphi[20] <= 1974; iphi[21] <= 2154; iphi[22] <= 2998; iphi[23] <= 1703; 
        iphi[24] <= 1919; iphi[25] <= 2266; iphi[26] <= 712; iphi[27] <= 1637; iphi[28] <= 56; iphi[29] <= 2186; iphi[30] <= 3296; iphi[31] <= 733; 
        iphi[32] <= 3289; iphi[33] <= 1292; iphi[34] <= 2877; iphi[35] <= 3281; iphi[36] <= 2882; iphi[37] <= 1455; iphi[38] <= 1274; iphi[39] <= 1461; 
        iphi[40] <= 1746; iphi[41] <= 863; iphi[42] <= 2419; iphi[43] <= 2761; iphi[44] <= 3033; iphi[45] <= 2237; iphi[46] <= 650; iphi[47] <= 2308; 
        iphi[48] <= 687; iphi[49] <= 780; iphi[50] <= 1438; iphi[51] <= 2156; iphi[52] <= 936; iphi[53] <= 394; iphi[54] <= 3253; iphi[55] <= 1789; 
        iphi[56] <= 3136; iphi[57] <= 2572; iphi[58] <= 1481; iphi[59] <= 1100; iphi[60] <= 1089; iphi[61] <= 2443; iphi[62] <= 1320; iphi[63] <= 641; 
        iphi[64] <= 1600; iphi[65] <= 1584; iphi[66] <= 1435; iphi[67] <= 1920; iphi[68] <= 1235; iphi[69] <= 1722; iphi[70] <= 2304; iphi[71] <= 1482; 
        iphi[72] <= 69; iphi[73] <= 2099; iphi[74] <= 3110; iphi[75] <= 2746; iphi[76] <= 1853; iphi[77] <= 403; iphi[78] <= 632; iphi[79] <= 892; 
        iphi[80] <= 2481; iphi[81] <= 2090; iphi[82] <= 2402; iphi[83] <= 314; iphi[84] <= 2508; iphi[85] <= 885; iphi[86] <= 3040; iphi[87] <= 1678; 
        iphi[88] <= 1062; iphi[89] <= 319; iphi[90] <= 682; iphi[91] <= 2606; iphi[92] <= 3046; iphi[93] <= 2150; iphi[94] <= 464; iphi[95] <= 992; 
        iphi[96] <= 2580; iphi[97] <= 3220; iphi[98] <= 2522; iphi[99] <= 3096; iphi[100] <= 535; iphi[101] <= 1029; iphi[102] <= 1052; iphi[103] <= 642; 
        iphi[104] <= 569; iphi[105] <= 2594; iphi[106] <= 2102; iphi[107] <= 17; iphi[108] <= 2447; iphi[109] <= 525; iphi[110] <= 1352; iphi[111] <= 939; 
        iphi[112] <= 630; iphi[113] <= 2954; iphi[114] <= 461; iphi[115] <= 756; iphi[116] <= 2879; iphi[117] <= 1219; iphi[118] <= 1573; iphi[119] <= 2789; 
        iphi[120] <= 797; iphi[121] <= 556; iphi[122] <= 2681; iphi[123] <= 2288; iphi[124] <= 1333; iphi[125] <= 554; iphi[126] <= 1414; iphi[127] <= 268;
    end
end



// for 2*N = 512, p = 1049089
else if (N == 256)
begin
    // phi = 841160 for 2*N = 512, p = 1049089
    phi[0] <= 1; phi[1] <= 841160; phi[2] <= 462262; phi[3] <= 907871; phi[4] <= 365501; phi[5] <= 896998; phi[6] <= 390723; phi[7] <= 907671; 
    phi[8] <= 1036830; phi[9] <= 764430; phi[10] <= 308920; phi[11] <= 194612; phi[12] <= 1031449; phi[13] <= 252416; phi[14] <= 267117; phi[15] <= 548234; 
    phi[16] <= 263354; phi[17] <= 364667; phi[18] <= 161010; phi[19] <= 928967; phi[20] <= 136426; phi[21] <= 444806; phi[22] <= 668555; phi[23] <= 712617; 
    phi[24] <= 639256; phi[25] <= 764565; phi[26] <= 563908; phi[27] <= 703731; phi[28] <= 850621; phi[29] <= 287868; phi[30] <= 716612; phi[31] <= 841389; 
    phi[32] <= 55526; phi[33] <= 807880; phi[34] <= 548338; phi[35] <= 669607; phi[36] <= 181821; phi[37] <= 161584; phi[38] <= 124778; phi[39] <= 55297; 
    phi[40] <= 165527; phi[41] <= 648329; phi[42] <= 486770; phi[43] <= 409212; phi[44] <= 370486; phi[45] <= 870865; phi[46] <= 967349; phi[47] <= 874660; 
    phi[48] <= 791722; phi[49] <= 33053; phi[50] <= 953891; phi[51] <= 213690; phi[52] <= 767496; phi[53] <= 644718; phi[54] <= 170665; phi[55] <= 281729; 
    phi[56] <= 451430; phi[57] <= 800716; phi[58] <= 445314; phi[59] <= 998612; phi[60] <= 545777; phi[61] <= 238564; phi[62] <= 750320; phi[63] <= 934266; 
    phi[64] <= 913194; phi[65] <= 348329; phi[66] <= 354830; phi[67] <= 884122; phi[68] <= 409399; phi[69] <= 304056; phi[70] <= 239472; phi[71] <= 786808; 
    phi[72] <= 1032562; phi[73] <= 676108; phi[74] <= 711113; phi[75] <= 735950; phi[76] <= 19435; phi[77] <= 1039802; phi[78] <= 712863; phi[79] <= 894083; 
    phi[80] <= 130316; phi[81] <= 444217; phi[82] <= 395323; phi[83] <= 154350; phi[84] <= 938627; phi[85] <= 547721; phi[86] <= 972942; phi[87] <= 318375; 
    phi[88] <= 218703; phi[89] <= 164796; phi[90] <= 526523; phi[91] <= 379906; phi[92] <= 828848; phi[93] <= 706950; phi[94] <= 845952; phi[95] <= 701044; 
    phi[96] <= 391407; phi[97] <= 311250; phi[98] <= 399160; phi[99] <= 687506; phi[100] <= 628422; phi[101] <= 24179; phi[102] <= 768286; phi[103] <= 38692; 
    phi[104] <= 274673; phi[105] <= 972032; phi[106] <= 697745; phi[107] <= 244972; phi[108] <= 684318; phi[109] <= 481826; phi[110] <= 302968; phi[111] <= 912089; 
    phi[112] <= 359383; phi[113] <= 461663; phi[114] <= 615751; phi[115] <= 430059; phi[116] <= 510371; phi[117] <= 715225; phi[118] <= 739437; phi[119] <= 940600; 
    phi[120] <= 497603; phi[121] <= 308438; phi[122] <= 752935; phi[123] <= 628033; phi[124] <= 128707; phi[125] <= 342587; phi[126] <= 419866; phi[127] <= 770888; 
    phi[128] <= 337358; phi[129] <= 824403; phi[130] <= 703946; phi[131] <= 207624; phi[132] <= 10743; phi[133] <= 778323; phi[134] <= 742429; phi[135] <= 926809; 
    phi[136] <= 886205; phi[137] <= 567049; phi[138] <= 132100; phi[139] <= 876387; phi[140] <= 486777; phi[141] <= 2798; phi[142] <= 459053; phi[143] <= 931428; 
    phi[144] <= 378589; phi[145] <= 859112; phi[146] <= 379516; phi[147] <= 92216; phi[148] <= 868078; phi[149] <= 319255; phi[150] <= 831758; phi[151] <= 957913; 
    phi[152] <= 47185; phi[153] <= 999552; phi[154] <= 223071; phi[155] <= 441998; phi[156] <= 190614; phi[157] <= 404014; phi[158] <= 623758; phi[159] <= 446799; 
    phi[160] <= 656213; phi[161] <= 900641; phi[162] <= 347634; phi[163] <= 91203; phi[164] <= 633266; phi[165] <= 990632; phi[166] <= 160399; phi[167] <= 1033817; 
    phi[168] <= 948374; phi[169] <= 703706; phi[170] <= 803401; phi[171] <= 271297; phi[172] <= 50706; phi[173] <= 96576; phi[174] <= 710534; phi[175] <= 481606; 
    phi[176] <= 936521; phi[177] <= 976082; phi[178] <= 1003762; phi[179] <= 831296; phi[180] <= 504923; phi[181] <= 496297; phi[182] <= 149661; phi[183] <= 264938; 
    phi[184] <= 419077; phi[185] <= 119896; phi[186] <= 695612; phi[187] <= 1041971; phi[188] <= 823132; phi[189] <= 611277; phi[190] <= 162462; phi[191] <= 104602; 
    phi[192] <= 972979; phi[193] <= 1017714; phi[194] <= 536973; phi[195] <= 185175; phi[196] <= 411903; phi[197] <= 1047073; phi[198] <= 598353; phi[199] <= 719929; 
    phi[200] <= 392369; phi[201] <= 659551; phi[202] <= 281468; phi[203] <= 168271; phi[204] <= 795569; phi[205] <= 585097; phi[206] <= 20861; phi[207] <= 376146; 
    phi[208] <= 21494; phi[209] <= 942303; phi[210] <= 986598; phi[211] <= 723874; phi[212] <= 500062; phi[213] <= 966459; phi[214] <= 242717; phi[215] <= 621430; 
    phi[216] <= 875482; phi[217] <= 875591; phi[218] <= 242199; phi[219] <= 272485; phi[220] <= 616058; phi[221] <= 590285; phi[222] <= 797790; phi[223] <= 373948; 
    phi[224] <= 695721; phi[225] <= 408579; phi[226] <= 853418; phi[227] <= 954850; phi[228] <= 136689; phi[229] <= 312107; phi[230] <= 549137; phi[231] <= 290398; 
    phi[232] <= 249831; phi[233] <= 630014; phi[234] <= 513335; phi[235] <= 228912; phi[236] <= 773771; phi[237] <= 956959; phi[238] <= 133630; phi[239] <= 618984; 
    phi[240] <= 661651; phi[241] <= 51592; phi[242] <= 511146; phi[243] <= 80867; phi[244] <= 204049; phi[245] <= 601906; phi[246] <= 506848; phi[247] <= 984970; 
    phi[248] <= 376539; phi[249] <= 134339; phi[250] <= 69783; phi[251] <= 40552; phi[252] <= 640574; phi[253] <= 526372; phi[254] <= 304515; phi[255] <= 267160; 
    //phi[512] <= 1; 
    
    
    // iphi = 781929 for 2*N = 512, p = 1049089
    iphi[0] <= 1; iphi[1] <= 781929; iphi[2] <= 744574; iphi[3] <= 522717; iphi[4] <= 408515; iphi[5] <= 1008537; iphi[6] <= 979306; iphi[7] <= 914750; 
    iphi[8] <= 672550; iphi[9] <= 64119; iphi[10] <= 542241; iphi[11] <= 447183; iphi[12] <= 845040; iphi[13] <= 968222; iphi[14] <= 537943; iphi[15] <= 997497; 
    iphi[16] <= 387438; iphi[17] <= 430105; iphi[18] <= 915459; iphi[19] <= 92130; iphi[20] <= 275318; iphi[21] <= 820177; iphi[22] <= 535754; iphi[23] <= 419075; 
    iphi[24] <= 799258; iphi[25] <= 758691; iphi[26] <= 499952; iphi[27] <= 736982; iphi[28] <= 912400; iphi[29] <= 94239; iphi[30] <= 195671; iphi[31] <= 640510; 
    iphi[32] <= 353368; iphi[33] <= 675141; iphi[34] <= 251299; iphi[35] <= 458804; iphi[36] <= 433031; iphi[37] <= 776604; iphi[38] <= 806890; iphi[39] <= 173498; 
    iphi[40] <= 173607; iphi[41] <= 427659; iphi[42] <= 806372; iphi[43] <= 82630; iphi[44] <= 549027; iphi[45] <= 325215; iphi[46] <= 62491; iphi[47] <= 106786; 
    iphi[48] <= 1027595; iphi[49] <= 672943; iphi[50] <= 1028228; iphi[51] <= 463992; iphi[52] <= 253520; iphi[53] <= 880818; iphi[54] <= 767621; iphi[55] <= 389538; 
    iphi[56] <= 656720; iphi[57] <= 329160; iphi[58] <= 450736; iphi[59] <= 2016; iphi[60] <= 637186; iphi[61] <= 863914; iphi[62] <= 512116; iphi[63] <= 31375; 
    iphi[64] <= 76110; iphi[65] <= 944487; iphi[66] <= 886627; iphi[67] <= 437812; iphi[68] <= 225957; iphi[69] <= 7118; iphi[70] <= 353477; iphi[71] <= 929193; 
    iphi[72] <= 630012; iphi[73] <= 784151; iphi[74] <= 899428; iphi[75] <= 552792; iphi[76] <= 544166; iphi[77] <= 217793; iphi[78] <= 45327; iphi[79] <= 73007; 
    iphi[80] <= 112568; iphi[81] <= 567483; iphi[82] <= 338555; iphi[83] <= 952513; iphi[84] <= 998383; iphi[85] <= 777792; iphi[86] <= 245688; iphi[87] <= 345383; 
    iphi[88] <= 100715; iphi[89] <= 15272; iphi[90] <= 888690; iphi[91] <= 58457; iphi[92] <= 415823; iphi[93] <= 957886; iphi[94] <= 701455; iphi[95] <= 148448; 
    iphi[96] <= 392876; iphi[97] <= 602290; iphi[98] <= 425331; iphi[99] <= 645075; iphi[100] <= 858475; iphi[101] <= 607091; iphi[102] <= 826018; iphi[103] <= 49537; 
    iphi[104] <= 1001904; iphi[105] <= 91176; iphi[106] <= 217331; iphi[107] <= 729834; iphi[108] <= 181011; iphi[109] <= 956873; iphi[110] <= 669573; iphi[111] <= 189977; 
    iphi[112] <= 670500; iphi[113] <= 117661; iphi[114] <= 590036; iphi[115] <= 1046291; iphi[116] <= 562312; iphi[117] <= 172702; iphi[118] <= 916989; iphi[119] <= 482040; 
    iphi[120] <= 162884; iphi[121] <= 122280; iphi[122] <= 306660; iphi[123] <= 270766; iphi[124] <= 1038346; iphi[125] <= 841465; iphi[126] <= 345143; iphi[127] <= 224686; 
    iphi[128] <= 711731; iphi[129] <= 278201; iphi[130] <= 629223; iphi[131] <= 706502; iphi[132] <= 920382; iphi[133] <= 421056; iphi[134] <= 296154; iphi[135] <= 740651; 
    iphi[136] <= 551486; iphi[137] <= 108489; iphi[138] <= 309652; iphi[139] <= 333864; iphi[140] <= 538718; iphi[141] <= 619030; iphi[142] <= 433338; iphi[143] <= 587426; 
    iphi[144] <= 689706; iphi[145] <= 137000; iphi[146] <= 746121; iphi[147] <= 567263; iphi[148] <= 364771; iphi[149] <= 804117; iphi[150] <= 351344; iphi[151] <= 77057; 
    iphi[152] <= 774416; iphi[153] <= 1010397; iphi[154] <= 280803; iphi[155] <= 1024910; iphi[156] <= 420667; iphi[157] <= 361583; iphi[158] <= 649929; iphi[159] <= 737839; 
    iphi[160] <= 657682; iphi[161] <= 348045; iphi[162] <= 203137; iphi[163] <= 342139; iphi[164] <= 220241; iphi[165] <= 669183; iphi[166] <= 522566; iphi[167] <= 884293; 
    iphi[168] <= 830386; iphi[169] <= 730714; iphi[170] <= 76147; iphi[171] <= 501368; iphi[172] <= 110462; iphi[173] <= 894739; iphi[174] <= 653766; iphi[175] <= 604872; 
    iphi[176] <= 918773; iphi[177] <= 155006; iphi[178] <= 336226; iphi[179] <= 9287; iphi[180] <= 1029654; iphi[181] <= 313139; iphi[182] <= 337976; iphi[183] <= 372981; 
    iphi[184] <= 16527; iphi[185] <= 262281; iphi[186] <= 809617; iphi[187] <= 745033; iphi[188] <= 639690; iphi[189] <= 164967; iphi[190] <= 694259; iphi[191] <= 700760; 
    iphi[192] <= 135895; iphi[193] <= 114823; iphi[194] <= 298769; iphi[195] <= 810525; iphi[196] <= 503312; iphi[197] <= 50477; iphi[198] <= 603775; iphi[199] <= 248373; 
    iphi[200] <= 597659; iphi[201] <= 767360; iphi[202] <= 878424; iphi[203] <= 404371; iphi[204] <= 281593; iphi[205] <= 835399; iphi[206] <= 95198; iphi[207] <= 1016036; 
    iphi[208] <= 257367; iphi[209] <= 174429; iphi[210] <= 81740; iphi[211] <= 178224; iphi[212] <= 678603; iphi[213] <= 639877; iphi[214] <= 562319; iphi[215] <= 400760; 
    iphi[216] <= 883562; iphi[217] <= 993792; iphi[218] <= 924311; iphi[219] <= 887505; iphi[220] <= 867268; iphi[221] <= 379482; iphi[222] <= 500751; iphi[223] <= 241209; 
    iphi[224] <= 993563; iphi[225] <= 207700; iphi[226] <= 332477; iphi[227] <= 761221; iphi[228] <= 198468; iphi[229] <= 345358; iphi[230] <= 485181; iphi[231] <= 284524; 
    iphi[232] <= 409833; iphi[233] <= 336472; iphi[234] <= 380534; iphi[235] <= 604283; iphi[236] <= 912663; iphi[237] <= 120122; iphi[238] <= 888079; iphi[239] <= 684422; 
    iphi[240] <= 785735; iphi[241] <= 500855; iphi[242] <= 781972; iphi[243] <= 796673; iphi[244] <= 17640; iphi[245] <= 854477; iphi[246] <= 740169; iphi[247] <= 284659; 
    iphi[248] <= 12259; iphi[249] <= 141418; iphi[250] <= 658366; iphi[251] <= 152091; iphi[252] <= 683588; iphi[253] <= 141218; iphi[254] <= 586827; iphi[255] <= 207929; 
    //iphi[512] <= 1;
end


